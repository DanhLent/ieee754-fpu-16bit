module Add_SubUnit_ver(
    input wire [15:0] Ain,
    input wire [15:0] Bin,
	 input wire Select,   // 0: Add, 1: Sub
	 input wire CLK,
	 input wire Start,
    input wire Reset,
	 output reg [15:0] Out,
    output reg Done
);

    // ============================================================
    // STAGE 1: DECODE & ALIGNMENT
    // ============================================================
    reg [4:0]  s1_exp_max;
    reg [11:0] s1_man_l, s1_man_s_shifted;
    reg        s1_sign_l, s1_real_op, s1_start;

    wire sign_a = Ain[15];
    wire sign_b = Bin[15];
    wire [4:0] exp_a = Ain[14:10];
    wire [4:0] exp_b = Bin[14:10];
    
    wire [10:0] man_a = (exp_a == 5'd0) ? {1'b0, Ain[9:0]} : {1'b1, Ain[9:0]};
    wire [10:0] man_b = (exp_b == 5'd0) ? {1'b0, Bin[9:0]} : {1'b1, Bin[9:0]};

    wire a_gt_b = (exp_a > exp_b) || (exp_a == exp_b && man_a > man_b);
    wire [4:0] exp_diff = a_gt_b ? (exp_a - exp_b) : (exp_b - exp_a);
    wire actual_sub = sign_a ^ sign_b ^ Select;

    always @(posedge CLK or posedge Reset) begin
        if (Reset) begin
            s1_start <= 1'b0;
            s1_exp_max <= 5'd0;
            s1_sign_l  <= 1'b0;
            s1_real_op <= 1'b0;
            s1_man_l   <= 12'd0;
            s1_man_s_shifted <= 12'd0;
        end else begin
            s1_start <= Start;
            s1_exp_max <= a_gt_b ? exp_a : exp_b;
            s1_sign_l  <= a_gt_b ? sign_a : (Select ? ~sign_b : sign_b);
            s1_real_op <= actual_sub;
            s1_man_l   <= a_gt_b ? {man_a, 1'b0} : {man_b, 1'b0};
            s1_man_s_shifted <= a_gt_b ? ({man_b, 1'b0} >> exp_diff) : ({man_a, 1'b0} >> exp_diff);
        end
    end

    // ============================================================
    // STAGE 2: ARITHMETIC (ADD/SUB)
    // ============================================================
    reg [12:0] s2_sum; // Sử dụng 13 bit để kiểm tra carry out dễ hơn
    reg [4:0]  s2_exp_max;
    reg        s2_sign_l, s2_real_op, s2_start;

    always @(posedge CLK or posedge Reset) begin
        if (Reset) begin
            s2_start <= 1'b0;
            s2_exp_max <= 5'd0;
            s2_sign_l  <= 1'b0;
            s2_real_op <= 1'b0;
            s2_sum <= 13'd0;
        end else begin
            s2_start <= s1_start;
            s2_exp_max <= s1_exp_max;
            s2_sign_l  <= s1_sign_l;
            s2_real_op <= s1_real_op;
            if (s1_real_op)
                s2_sum <= {1'b0, s1_man_l} - {1'b0, s1_man_s_shifted};
            else
                s2_sum <= {1'b0, s1_man_l} + {1'b0, s1_man_s_shifted};
        end
    end

    // ============================================================
    // STAGE 3: NORMALIZATION & PACKING
    // ============================================================
    reg [3:0] l_zeros;
    
    // Tìm vị trí bit 1 đầu tiên
    always @(*) begin
        if      (s2_sum[12]) l_zeros = 4'd0; 
        else if (s2_sum[11]) l_zeros = 4'd0; 
        else if (s2_sum[10]) l_zeros = 4'd1;
        else if (s2_sum[9])  l_zeros = 4'd2;
        else if (s2_sum[8])  l_zeros = 4'd3;
        else if (s2_sum[7])  l_zeros = 4'd4;
        else if (s2_sum[6])  l_zeros = 4'd5;
        else if (s2_sum[5])  l_zeros = 4'd6;
        else if (s2_sum[4])  l_zeros = 4'd7;
        else if (s2_sum[3])  l_zeros = 4'd8;
        else if (s2_sum[2])  l_zeros = 4'd9;
        else if (s2_sum[1])  l_zeros = 4'd10;
        else if (s2_sum[0])  l_zeros = 4'd11;
        else                 l_zeros = 4'd12;
    end

    // Tính toán các thành phần trung gian để tránh lỗi cú pháp trong dấu {}
    wire [4:0] final_exp_norm = s2_exp_max - l_zeros;
    wire [11:0] shifted_man    = s2_sum[11:0] << l_zeros;
    wire [9:0]  final_man_norm = shifted_man[10:1]; // Bỏ bit ẩn sau khi dịch

    always @(posedge CLK or posedge Reset) begin
        if (Reset) begin
            Done <= 1'b0;
            Out  <= 16'h0000;
        end else begin
            Done <= s2_start;
            if (s2_sum == 13'd0) begin
                Out <= 16'h0000;
            end else if (s2_sum[12]) begin
                // Trường hợp tràn (Cout)
                Out <= {s2_sign_l, (s2_exp_max + 5'd1), s2_sum[11:2]};
            end else if (s2_exp_max < l_zeros) begin
                // Trường hợp Underflow
                Out <= 16'h0000;
            end else begin
                // Trường hợp chuẩn hóa thông thường
                Out <= {s2_sign_l, final_exp_norm, final_man_norm};
            end
        end
    end

endmodule