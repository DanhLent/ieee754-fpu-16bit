module Add_SubUni1(
    input wire [15:0] Ain,
    input wire [15:0] Bin,
    input wire Select,
    input wire CLK,
    input wire Start,
    output reg [15:0] Out,
    output reg Done
);

    reg [4:0]  s1_exp_max;
    reg [11:0] s1_man_l, s1_man_s_shifted;
    reg        s1_sign_l, s1_real_op, s1_start;

    wire sign_a = Ain[15];
    wire sign_b = Bin[15];
    wire [4:0] exp_a = Ain[14:10];
    wire [4:0] exp_b = Bin[14:10];
    
    wire [10:0] man_a = (exp_a == 5'd0) ? {1'b0, Ain[9:0]} : {1'b1, Ain[9:0]};
    wire [10:0] man_b = (exp_b == 5'd0) ? {1'b0, Bin[9:0]} : {1'b1, Bin[9:0]};

    wire a_gt_b = (exp_a > exp_b) || (exp_a == exp_b && man_a > man_b);
    wire [4:0] exp_diff = a_gt_b ? (exp_a - exp_b) : (exp_b - exp_a);
    wire actual_sub = sign_a ^ sign_b ^ Select;

    always @(posedge CLK) begin
        s1_start <= Start;
        s1_exp_max <= a_gt_b ? exp_a : exp_b;
        s1_sign_l  <= a_gt_b ? sign_a : (Select ? ~sign_b : sign_b);
        s1_real_op <= actual_sub;
        s1_man_l   <= a_gt_b ? {man_a, 1'b0} : {man_b, 1'b0};
        s1_man_s_shifted <= a_gt_b ? ({man_b, 1'b0} >> exp_diff) : ({man_a, 1'b0} >> exp_diff);
    end

    reg [12:0] s2_sum;
    reg [4:0]  s2_exp_max;
    reg        s2_sign_l, s2_real_op, s2_start;

    always @(posedge CLK) begin
        s2_start <= s1_start;
        s2_exp_max <= s1_exp_max;
        s2_sign_l  <= s1_sign_l;
        s2_real_op <= s1_real_op;
        if (s1_real_op)
            s2_sum <= {1'b0, s1_man_l} - {1'b0, s1_man_s_shifted};
        else
            s2_sum <= {1'b0, s1_man_l} + {1'b0, s1_man_s_shifted};
    end

    reg [3:0] l_zeros;
    
    always @(*) begin
        if      (s2_sum[12]) l_zeros = 4'd0;
        else if (s2_sum[11]) l_zeros = 4'd0; 
        else if (s2_sum[10]) l_zeros = 4'd1;
        else if (s2_sum[9])  l_zeros = 4'd2;
        else if (s2_sum[8])  l_zeros = 4'd3;
        else if (s2_sum[7])  l_zeros = 4'd4;
        else if (s2_sum[6])  l_zeros = 4'd5;
        else if (s2_sum[5])  l_zeros = 4'd6;
        else if (s2_sum[4])  l_zeros = 4'd7;
        else if (s2_sum[3])  l_zeros = 4'd8;
        else if (s2_sum[2])  l_zeros = 4'd9;
        else if (s2_sum[1])  l_zeros = 4'd10;
        else if (s2_sum[0])  l_zeros = 4'd11;
        else                 l_zeros = 4'd12;
    end

    wire [4:0] final_exp_norm = s2_exp_max - l_zeros;
    wire [11:0] shifted_man    = s2_sum[11:0] << l_zeros;
    wire [9:0]  final_man_norm = shifted_man[10:1]; 

    always @(posedge CLK) begin
        Done <= s2_start;
        if (s2_sum == 13'd0) begin
            Out <= 16'h0000;
        end else if (s2_sum[12]) begin
            Out <= {s2_sign_l, (s2_exp_max + 5'd1), s2_sum[11:2]};
        end else if (s2_exp_max < l_zeros) begin
            Out <= 16'h0000;
        end else begin
            Out <= {s2_sign_l, final_exp_norm, final_man_norm};
        end
    end

endmodule